`define CYCLE_PCI       2'b00
`define CYCLE_PCR       2'b10
`define CYCLE_PCC       2'b01
`define CYCLE_PCW       2'b11

`define REG_A           3'b000
`define REG_B           3'b001
`define REG_C           3'b010
`define REG_D           3'b011
`define REG_E           3'b100
`define REG_H           3'b101
`define REG_L           3'b110
`define REG_M           3'b111

`define STATE_T1        3'b010
`define STATE_T1I       3'b110
`define STATE_T2        3'b100
`define STATE_WAIT      3'b000
`define STATE_T3        3'b001
`define STATE_STOPPED   3'b011
`define STATE_T4        3'b111
`define STATE_T5        3'b101
